library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package Types is
    type sound is (blaster, victory, game_over);
end Types;

package body Types is

end Types;
